//Hayden Prater
//November 21, 2022
//Memory Load/Store

module MemLoadStore ();
    // Fill In code

endmodule